module ParityGenerator(
input x,y,z,
output result);
xor (result,x,y,z);  
endmodule